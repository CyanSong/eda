title
*netlist example 1
r1 1 0 5
L3 2 0 4m

cap2 1 0 3
v3 1 2 ac 1
r4 2 0 8
.end