title
*netlist example 1
r1 1 0 5
g2 1 0 1 2 2
h2 1 0 v3 4
v3 1 2 6
r4 2 0 8
is 0 2 10
.end