title

*netlist example 1

r1 0 1 1
c1 1 2 1
v1 2 0 1
.tran .2 5 0
.plot tran   v(1)



.end